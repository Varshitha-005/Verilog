module test;
 initial begin
    $display("Hello Verilog from VS Code");
    $finish;
 end
endmodule